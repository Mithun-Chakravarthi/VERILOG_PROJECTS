module dct_test_final;

    reg signed [0:511] A; 
    reg clk;              
    reg reset;          
    wire signed [103:0] D; 
    integer i, j;

    dct_final dat (
        .A(A),
        .clk(clk),
        .reset(reset),
        .D(D));

    always #5 clk = ~clk; 

    initial begin
        clk = 0;
        reset = 1; 
        A = 512'd0; 

        #10;
        reset = 0; 

    // Initialize A with specified values
/*A ={-8'd102, -8'd16, -8'd19, -8'd12, -8'd12, -8'd27, -8'd51, -8'd47,  // Row 1
     -8'd106, -8'd24, -8'd12, -8'd19, -8'd12, -8'd20, -8'd39, -8'd51,  // Row 2
     -8'd24, 8'd27, 8'd8, 8'd39, 8'd35, 8'd34, 8'd24, -8'd44,  // Row 3
     -8'd40, 8'd17, 8'd28, 8'd32, 8'd24, 8'd27, 8'd8, -8'd32,  // Row 4
     -8'd34, 8'd20, 8'd28, 8'd20, 8'd12, 8'd8, 8'd19, -8'd34,  // Row 5
     -8'd19, 8'd39, 8'd12, 8'd27, 8'd27, 8'd12, 8'd8, -8'd34,  // Row 6
     -8'd80, 8'd28, -8'd5, 8'd39, 8'd34, 8'd16, 8'd12, -8'd19,  // Row 7
     -8'd120, -8'd27, -8'd8, -8'd27, -8'd24, -8'd19, -8'd19, -8'd8};   // Row 8*/
A = {8'd26, 8'd112, 8'd109, 8'd116, 8'd116, 8'd101, 8'd77, 8'd81, 
     8'd22, 8'd104, 8'd116, 8'd109, 8'd116, 8'd108, 8'd89, 8'd77, 
     8'd104, 8'd155, 8'd136, 8'd167, 8'd163, 8'd162, 8'd152, 8'd84, 
     8'd88, 8'd145, 8'd156, 8'd160, 8'd152, 8'd155, 8'd136, 8'd96, 
     8'd94, 8'd148, 8'd156, 8'd148, 8'd140, 8'd136, 8'd147, 8'd94, 
     8'd109, 8'd167, 8'd140, 8'd155, 8'd155, 8'd140, 8'd136, 8'd94, 
     8'd48, 8'd156, 8'd123, 8'd167, 8'd162, 8'd144, 8'd140, 8'd109, 
     8'd8, 8'd101, 8'd120, 8'd101, 8'd104, 8'd109, 8'd109, 8'd120};


 /*
A = {-8'd76, -8'd73, -8'd67, -8'd62, -8'd58, -8'd67, -8'd64, -8'd55,  
     -8'd65, -8'd69, -8'd73, -8'd38, -8'd19, -8'd43, -8'd59, -8'd56, 
     -8'd66, -8'd69, -8'd60, -8'd15, 8'd16, -8'd24, -8'd62, -8'd55,  
     -8'd65, -8'd70, -8'd57, -8'd6, 8'd26, -8'd22, -8'd58, -8'd59,  
     -8'd61, -8'd67, -8'd60, -8'd24, -8'd2, -8'd40, -8'd60, -8'd58, 
     -8'd49, -8'd63, -8'd68, -8'd58, -8'd51, -8'd60, -8'd70, -8'd53,  
     -8'd43, -8'd57, -8'd64, -8'd69, -8'd73, -8'd67, -8'd63, -8'd45,  
     -8'd41, -8'd49, -8'd59, -8'd60, -8'd63, -8'd52, -8'd50, -8'd34};

A = {8'd52, 8'd55, 8'd61, 8'd66, 8'd70, 8'd61, 8'd64, 8'd73, 8'd63, 
     8'd59,8'd55, 8'd90, 8'd109, 8'd85, 8'd69, 8'd72, 8'd62, 8'd59, 8'd68, 8'd113, 
     8'd144, 8'd104, 8'd66, 8'd73, 8'd63, 8'd58, 8'd71, 8'd122, 8'd154, 8'd106, 
     8'd70, 8'd69, 8'd67, 8'd61, 8'd68, 8'd104, 8'd126, 8'd88, 8'd68, 8'd70, 
     8'd79, 8'd65, 8'd60, 8'd70, 8'd77, 8'd68, 8'd58, 8'd75, 8'd85, 8'd71, 
     8'd64, 8'd59, 8'd55, 8'd61, 8'd65, 8'd83, 8'd87, 8'd79, 8'd69, 8'd68, 
     8'd65, 8'd76, 8'd78, 8'd94};
*/
/*
A = {8'd52, 8'd55, 8'd61, 8'd66, 8'd70, 8'd61, 8'd64, 8'd73,    // Row 1
     8'd63, 8'd59, 8'd55, 8'd90, 8'd109, 8'd85, 8'd69, 8'd72,   // Row 2
     8'd62, 8'd59, 8'd68, 8'd113, 8'd144, 8'd104, 8'd66, 8'd73, // Row 3
     8'd63, 8'd58, 8'd71, 8'd122, 8'd154, 8'd106, 8'd70, 8'd69, // Row 4
     8'd67, 8'd61, 8'd68, 8'd104, 8'd126, 8'd88, 8'd68, 8'd70,  // Row 5
     8'd79, 8'd65, 8'd60, 8'd70, 8'd77, 8'd68, 8'd58, 8'd75,    // Row 6
     8'd85, 8'd71, 8'd64, 8'd59, 8'd55, 8'd61, 8'd65, 8'd83,    // Row 7
     8'd87, 8'd79, 8'd69, 8'd68, 8'd65, 8'd76, 8'd78, 8'd94};   // Row 8
*/
/*
A = {8'd39, 8'd43, 8'd46, 8'd39, 8'd39, 8'd54, 8'd78, 8'd74,  // Row 1
     8'd43, 8'd51, 8'd39, 8'd46, 8'd39, 8'd47, 8'd66, 8'd78,  // Row 2
     8'd51, 8'd54, 8'd35, 8'd66, 8'd62, 8'd61, 8'd51, 8'd71,  // Row 3
     8'd67, 8'd44, 8'd55, 8'd59, 8'd51, 8'd54, 8'd35, 8'd59,  // Row 4
     8'd61, 8'd47, 8'd55, 8'd47, 8'd39, 8'd35, 8'd46, 8'd61,  // Row 5
     8'd46, 8'd66, 8'd39, 8'd54, 8'd54, 8'd39, 8'd35, 8'd61,  // Row 6
     8'd35, 8'd55, 8'd22, 8'd66, 8'd61, 8'd43, 8'd39, 8'd46,  // Row 7
     8'd47, 8'd54, 8'd35, 8'd54, 8'd51, 8'd46, 8'd46, 8'd35};  // Row 8
*/
        #200;
        for (i = 0; i <= 7; i = i + 1) begin
            for (j = 0; j <= 7; j = j + 1) begin
                $display("matD[%0d][%0d] = %d", i, j, dat.matD[i][j]);
            end
        end
        
        #200;
        $finish; 
    end

endmodule

